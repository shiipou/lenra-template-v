module listeners

import x.json2 { Any }
import src.data { Api, Counter, SavedCounter }

pub fn on_session_start(props map[string]Any, event map[string]Any, api Api) ! {
}
